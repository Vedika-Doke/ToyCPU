// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Wed Nov 19 10:31:30 2025"

module C16dmuxer(
	DMUX_SEL
);


input wire	[4:0] DMUX_SEL;

wire	[15:0] DMUXOUT;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_79;




assign	SYNTHESIZED_WIRE_78 =  ~SYNTHESIZED_WIRE_72;

assign	SYNTHESIZED_WIRE_76 =  ~SYNTHESIZED_WIRE_73;

assign	SYNTHESIZED_WIRE_75 =  ~SYNTHESIZED_WIRE_74;



assign	SYNTHESIZED_WIRE_74 =  ~SYNTHESIZED_WIRE_11;

assign	SYNTHESIZED_WIRE_12 = ;

assign	SYNTHESIZED_WIRE_73 =  ~SYNTHESIZED_WIRE_12;

assign	SYNTHESIZED_WIRE_13 = ;

assign	SYNTHESIZED_WIRE_72 =  ~SYNTHESIZED_WIRE_13;


assign	SYNTHESIZED_WIRE_22 = ;


assign	SYNTHESIZED_WIRE_77 =  ~SYNTHESIZED_WIRE_22;













assign	SYNTHESIZED_WIRE_79 =  ~SYNTHESIZED_WIRE_77;

assign	SYNTHESIZED_WIRE_11 = ;


endmodule
