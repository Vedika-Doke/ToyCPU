// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Wed Nov 19 10:28:49 2025"

module Control_FSM(
	NOOP,
	INPUT_DATAC,
	INPUT_DATACF,
	INPUT_DATAD,
	INPUT_DATADF,
	MOVE,
	ADD,
	ADDI,
	SUB,
	SUBI,
	LOAD,
	LOADF,
	STORE,
	STOREF,
	SHIFTL,
	SHIFTR,
	CMP,
	ZERO_FLAG,
	JUMP,
	BRE/BRZ,
	BRNE/BRNZ,
	BRG,
	CARRY_FLAG,
	OVERFLOW_FLAG,
	NEGATIVE_FLAG,
	BRGE,
	LOADI/LOADP,
	X,
	Y,
	IMEM_WRITE_ENABLE,
	ALU_SOURCE_MUX,
	ALU_SELECT1,
	DMEM_WRITE_ENABLE,
	REG_WRITEBACK_MUX,
	ALU_SELECT0,
	PC_WRITE_ENABLE,
	PC_MUX,
	DMEM_INPUT_MUX,
	ALU_RESULT_MUX,
	FLAGS_WRITE_ENABLE,
	REG_WRITE_ENABLE,
	REG_PORT0_SELECT,
	REG_PORT1_SELECT,
	REG_WRITE_SELECT
);


input wire	NOOP;
input wire	INPUT_DATAC;
input wire	INPUT_DATACF;
input wire	INPUT_DATAD;
input wire	INPUT_DATADF;
input wire	MOVE;
input wire	ADD;
input wire	ADDI;
input wire	SUB;
input wire	SUBI;
input wire	LOAD;
input wire	LOADF;
input wire	STORE;
input wire	STOREF;
input wire	SHIFTL;
input wire	SHIFTR;
input wire	CMP;
input wire	ZERO_FLAG;
input wire	JUMP;
input wire	BRE/BRZ;
input wire	BRNE/BRNZ;
input wire	BRG;
input wire	CARRY_FLAG;
input wire	OVERFLOW_FLAG;
input wire	NEGATIVE_FLAG;
input wire	BRGE;
input wire	LOADI/LOADP;
input wire	[1:0] X;
input wire	[1:0] Y;
output wire	IMEM_WRITE_ENABLE;
output wire	ALU_SOURCE_MUX;
output wire	ALU_SELECT1;
output wire	DMEM_WRITE_ENABLE;
output wire	REG_WRITEBACK_MUX;
output wire	ALU_SELECT0;
output wire	PC_WRITE_ENABLE;
output wire	PC_MUX;
output wire	DMEM_INPUT_MUX;
output wire	ALU_RESULT_MUX;
output wire	FLAGS_WRITE_ENABLE;
output wire	REG_WRITE_ENABLE;
output wire	[1:0] REG_PORT0_SELECT;
output wire	[1:0] REG_PORT1_SELECT;
output wire	[1:0] REG_WRITE_SELECT;

wire	[1:0] REG_PORT0_SELECT_ALTERA_SYNTHESIZED;
wire	[1:0] REG_PORT1_SELECT_ALTERA_SYNTHESIZED;
wire	[1:0] REG_WRITE_SELECT_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;

assign	PC_WRITE_ENABLE = 1;
assign	REG_WRITE_ENABLE = SYNTHESIZED_WIRE_49;




assign	IMEM_WRITE_ENABLE = INPUT_DATAC | INPUT_DATACF;

assign	SYNTHESIZED_WIRE_36 = BRE/BRZ & ZERO_FLAG;

assign	SYNTHESIZED_WIRE_39 = SYNTHESIZED_WIRE_43 & BRNE/BRNZ;

assign	SYNTHESIZED_WIRE_37 = BRG & SYNTHESIZED_WIRE_1;

assign	SYNTHESIZED_WIRE_38 = SYNTHESIZED_WIRE_44 & BRGE;

assign	SYNTHESIZED_WIRE_45 = SUB | CMP | ADD;

assign	SYNTHESIZED_WIRE_43 =  ~ZERO_FLAG;

assign	SYNTHESIZED_WIRE_44 = OVERFLOW_FLAG ~^ NEGATIVE_FLAG;

assign	SYNTHESIZED_WIRE_1 = SYNTHESIZED_WIRE_43 & SYNTHESIZED_WIRE_44;

assign	SYNTHESIZED_WIRE_5 = STOREF | STORE;

assign	SYNTHESIZED_WIRE_48 = SYNTHESIZED_WIRE_5 | SYNTHESIZED_WIRE_45;

assign	SYNTHESIZED_WIRE_13 = SUB | LOAD | SUBI | LOADF | SHIFTL | SHIFTR;

assign	SYNTHESIZED_WIRE_46 = LOADF | STOREF | MOVE;

assign	SYNTHESIZED_WIRE_32 = SHIFTR | CMP | SHIFTL;

assign	SYNTHESIZED_WIRE_9 = INPUT_DATADF | ADD | INPUT_DATACF;

assign	SYNTHESIZED_WIRE_7 = SUB | SUBI | ADDI;

assign	SYNTHESIZED_WIRE_8 = SHIFTR | CMP | SHIFTL;

assign	SYNTHESIZED_WIRE_11 = SYNTHESIZED_WIRE_7 | SYNTHESIZED_WIRE_8 | SYNTHESIZED_WIRE_9;


Block3	b2v_inst43(
	.i0(X[1]),
	.i1(Y[1]),
	.sel(SYNTHESIZED_WIRE_46),
	.mxout(SYNTHESIZED_WIRE_15));

assign	SYNTHESIZED_WIRE_47 = SYNTHESIZED_WIRE_11 | SYNTHESIZED_WIRE_46;

assign	SYNTHESIZED_WIRE_29 = STOREF | CMP | LOADF;

assign	ALU_SELECT0 = SUB | SHIFTR | CMP | SUBI;

assign	SYNTHESIZED_WIRE_14 = MOVE | ADD | ADDI | LOADI/LOADP;

assign	SYNTHESIZED_WIRE_49 = SYNTHESIZED_WIRE_13 | SYNTHESIZED_WIRE_14;

assign	REG_PORT0_SELECT_ALTERA_SYNTHESIZED[1] = SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_47;


Block3	b2v_inst50(
	.i0(X[0]),
	.i1(Y[0]),
	.sel(SYNTHESIZED_WIRE_46),
	.mxout(SYNTHESIZED_WIRE_18));

assign	REG_PORT0_SELECT_ALTERA_SYNTHESIZED[0] = SYNTHESIZED_WIRE_18 & SYNTHESIZED_WIRE_47;

assign	REG_PORT1_SELECT_ALTERA_SYNTHESIZED[1] = SYNTHESIZED_WIRE_20 & SYNTHESIZED_WIRE_48;

assign	REG_PORT1_SELECT_ALTERA_SYNTHESIZED[0] = SYNTHESIZED_WIRE_22 & SYNTHESIZED_WIRE_48;

assign	REG_WRITE_SELECT_ALTERA_SYNTHESIZED[1] = X[1] & SYNTHESIZED_WIRE_49;

assign	REG_WRITE_SELECT_ALTERA_SYNTHESIZED[0] = X[0] & SYNTHESIZED_WIRE_49;

assign	SYNTHESIZED_WIRE_27 = INPUT_DATADF | MOVE | INPUT_DATACF;

assign	SYNTHESIZED_WIRE_26 = ADDI | LOADF | STOREF | SUBI;

assign	ALU_SOURCE_MUX = SYNTHESIZED_WIRE_26 | SYNTHESIZED_WIRE_27;

assign	SYNTHESIZED_WIRE_28 = ADD | SUB | SUBI | ADDI;

assign	SYNTHESIZED_WIRE_30 = INPUT_DATADF | MOVE | INPUT_DATACF;

assign	ALU_SELECT1 = SYNTHESIZED_WIRE_28 | SYNTHESIZED_WIRE_29 | SYNTHESIZED_WIRE_30;


Block3	b2v_inst64(
	.i0(X[1]),
	.i1(Y[1]),
	.sel(SYNTHESIZED_WIRE_45),
	.mxout(SYNTHESIZED_WIRE_20));

assign	SYNTHESIZED_WIRE_33 = ADD | SUB | SUBI | ADDI;

assign	FLAGS_WRITE_ENABLE = SYNTHESIZED_WIRE_32 | SYNTHESIZED_WIRE_33;

assign	SYNTHESIZED_WIRE_35 = INPUT_DATAD | LOADI/LOADP | INPUT_DATAC;

assign	SYNTHESIZED_WIRE_34 = STORE | LOAD;

assign	ALU_RESULT_MUX = SYNTHESIZED_WIRE_34 | SYNTHESIZED_WIRE_35;

assign	DMEM_INPUT_MUX = INPUT_DATADF | INPUT_DATAD;

assign	DMEM_WRITE_ENABLE = INPUT_DATAD | STORE | STOREF | INPUT_DATADF;

assign	REG_WRITEBACK_MUX = LOADF | LOAD;

assign	SYNTHESIZED_WIRE_41 = SYNTHESIZED_WIRE_36 | JUMP;

assign	SYNTHESIZED_WIRE_40 = SYNTHESIZED_WIRE_37 | SYNTHESIZED_WIRE_38 | SYNTHESIZED_WIRE_39;

assign	PC_MUX = SYNTHESIZED_WIRE_40 | SYNTHESIZED_WIRE_41;


Block3	b2v_inst76(
	.i0(X[0]),
	.i1(Y[0]),
	.sel(SYNTHESIZED_WIRE_45),
	.mxout(SYNTHESIZED_WIRE_22));

assign	REG_PORT0_SELECT = REG_PORT0_SELECT_ALTERA_SYNTHESIZED;
assign	REG_PORT1_SELECT = REG_PORT1_SELECT_ALTERA_SYNTHESIZED;
assign	REG_WRITE_SELECT = REG_WRITE_SELECT_ALTERA_SYNTHESIZED;

endmodule
